///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ZicsrM_mcause_cg = new();      ZicsrM_mcause_cg.set_inst_name("obj_ZicsrM_mcause");
    ZicsrM_mstatus_cg = new();     ZicsrM_mstatus_cg.set_inst_name("obj_ZicsrM_mstatus");
    ZicsrM_mprivinst_cg = new();   ZicsrM_mprivinst_cg.set_inst_name("obj_ZicsrM_mprivinst");
