///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ExceptionsVMZalrsc_cg = new();         ExceptionsVMZalrsc_cg.set_inst_name("obj_ExceptionsVMZalrsc");
