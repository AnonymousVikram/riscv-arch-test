///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Written: Vikram Krishna vkrishna@hmc.edu October 9 2025
//
// Copyright (C) 2025 Harvey Mudd College
//
// SPDX-License-Identifier: Apache-2.0
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ZicsrH_csr_access_cg = new();    ZicsrH_csr_access_cg.set_inst_name("obj_ZicsrH_csr_access");
    ZicsrH_csr_walk_cg = new();      ZicsrH_csr_walk_cg.set_inst_name("obj_ZicsrH_csr_walk");
    ZicsrH_replica_cg = new();        ZicsrH_replica_cg.set_inst_name("obj_ZicsrH_replica");
    ZicsrH_hstatus_vgein_cg = new();  ZicsrH_hstatus_vgein_cg.set_inst_name("obj_ZicsrH_hstatus_vgein");
    ZicsrH_vscause_cg = new();      ZicsrH_vscause_cg.set_inst_name("obj_ZicsrH_vscause");
    ZicsrH_vsstatus_cg = new();     ZicsrH_vsstatus_cg.set_inst_name("obj_ZicsrH_vsstatus");
    ZicsrH_tvm_cg = new();        ZicsrH_tvm_cg.set_inst_name("obj_ZicsrH_tvm");
    ZicsrH_mtval_cg = new();      ZicsrH_mtval_cg.set_inst_name("obj_ZicsrH_mtval");
    ZicsrH_hprivinst_cg = new();   ZicsrH_hprivinst_cg.set_inst_name("obj_ZicsrH_hprivinst");
